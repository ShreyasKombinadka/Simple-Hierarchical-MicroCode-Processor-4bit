module CPU4_tb ;
